`default_nettype none

module tt_um_kercrafter_leds_racer (
    input wire clk,
    input wire GREEN_BTN,
    input wire RED_BTN,
    input wire BLUE_BTN,
    input wire YELLOW_BTN,
    input wire FORCE_RESET,
    output wire LEDS_LINE,
    output wire TP_SCREEN_0,
    output wire TP_SCREEN_1,
    output wire TP_BLUE_RTP,
    output wire TP_RED_RTP,
    output wire TP_GREEN_RTP,
    output wire TP_YELLOW_RTP,
    output wire TP_UPDATE_FRAME
);

endmodule

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity end_screen is
  generic (
    max_pos : integer := 109
  );

  port (
    enable : in std_logic;

    red_pos : in integer range 0 to max_pos-1;
    blue_pos : in integer range 0 to max_pos-1;
    green_pos : in integer range 0 to max_pos-1;
    yellow_pos : in integer range 0 to max_pos-1;
    
    led_number : in integer range 0 to max_pos-1;

    i_red_intensity : in std_logic_vector(7 downto 0);
    i_blue_intensity : in std_logic_vector(7 downto 0);
    i_green_intensity : in std_logic_vector(7 downto 0);
  
    o_red_intensity : out std_logic_vector(7 downto 0);
    o_blue_intensity : out std_logic_vector(7 downto 0);
    o_green_intensity : out std_logic_vector(7 downto 0)
  );
end entity;


architecture beh of end_screen is
    signal red_intensity : std_logic_vector(7 downto 0);
    signal blue_intensity : std_logic_vector(7 downto 0);
    signal green_intensity : std_logic_vector(7 downto 0);
begin

  pipe_tri_bus: entity work.pipe_tri_bus
    port map(
      enable => enable,

      i_led_red_intensity => i_red_intensity,
      i_led_blue_intensity => i_blue_intensity,
      i_led_green_intensity => i_green_intensity,

      d_led_green_intensity => green_intensity,
      d_led_red_intensity => red_intensity,
      d_led_blue_intensity => blue_intensity,

      o_led_green_intensity => o_green_intensity,
      o_led_red_intensity => o_red_intensity,
      o_led_blue_intensity => o_blue_intensity
    );

  process(led_number, red_pos, blue_pos, green_pos, yellow_pos)
    procedure set_GRB (green_intensity_i: integer range 0 to 255; red_intensity_i: integer range 0 to 255; blue_intensity_i: integer range 0 to 255) is
    begin
      green_intensity <= std_logic_vector(to_unsigned(green_intensity_i, 8));
      red_intensity <= std_logic_vector(to_unsigned(red_intensity_i, 8));
      blue_intensity <= std_logic_vector(to_unsigned(blue_intensity_i, 8));
    end procedure;
    
    procedure set_LED_white is
    begin
      set_GRB(5, 5, 5);
    end procedure;
    
    procedure set_LED_off is
    begin
      set_GRB(0, 0, 0);
    end procedure;
    
    procedure set_LED_green is
    begin
      set_GRB(5, 0, 0);
    end procedure;

    procedure set_LED_red is
    begin
      set_GRB(0, 5, 0);
    end procedure;
    
    procedure set_LED_blue is
    begin
      set_GRB(0, 0, 5);
    end procedure;

    procedure set_LED_yellow is
    begin
      set_GRB(5, 5, 0);
    end procedure;
  begin
    if green_pos = max_pos-1 then
      set_LED_green;
    elsif red_pos = max_pos-1 then
      set_LED_red;
    elsif blue_pos = max_pos-1 then
      set_LED_blue;
    elsif yellow_pos = max_pos-1 then
      set_LED_yellow;
    else
      set_LED_off;
    end if;
  end process;

end architecture;
